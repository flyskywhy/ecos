# ====================================================================
#
#      spi_microblaze.cdl
#
#      Microblaze SPI driver configuration data 
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2009 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Savin Zlobec <savin@elatec.si> 
# Contributors:   Li Zheng
# Date:           2004-08-25
# Description:    Ref to packages/devs/spi/arm/lpc2xxx/current/cdl/spi_lpc2xxx.cdl
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_SPI_MICROBLAZE {
    parent        CYGPKG_IO_SPI
    active_if     CYGPKG_IO_SPI
    display       "Microblaze SPI driver"
    description   "Microblaze SPI driver"
    hardware
    active_if     CYGPKG_HAL_MICROBLAZE
    requires      CYGPKG_HAL_MICROBLAZE_GENERIC
    
    active_if     MON_SPI_0
    
    include_dir   cyg/io
    compile       -library=libextras.a spi_microblaze.cxx spi_devices.c src/xspi.c src/xspi_g.c src/xspi_options.c \
                  src/xspi_selftest.c src/xspi_sinit.c src/xspi_stats.c src/xil_io.c

    cdl_component CYGPKG_DEVS_SPI_MICROBLAZE_BUS0 {
        active_if     MON_SPI_0
        display       "Enable SPI interface 0"
        flavor        bool
        default_value 1
        description   "Enable this component to get support for SPI interface 0."

        cdl_option CYGNUM_IO_SPI_MICROBLAZE_BUS0_INTPRIO {
            display       "Interrupt priority of the SPI bus 0 ISR"
            flavor        data
            legal_values  0 to 15
            default_value 12
            requires      { is_active(CYGNUM_IO_SPI_MICROBLAZE_BUS1_INTPRIO)
                             implies (CYGNUM_IO_SPI_MICROBLAZE_BUS0_INTPRIO !=
                             CYGNUM_IO_SPI_MICROBLAZE_BUS1_INTPRIO)
            }
            description "
                This option specifies the interrupt priority of the ISR of
                the SPI bus 0 interrupt in the VIC. Slot 0 has the highest
                priority and slot 15 the lowest."
        }
    }

    cdl_component CYGPKG_DEVS_SPI_MICROBLAZE_BUS1 {
        active_if     MON_SPI_1
        display       "Enable SPI interface 1"
        flavor        bool
        default_value 1
        description   "Enable this component to get support for SPI interface 1."

        cdl_option CYGNUM_IO_SPI_MICROBLAZE_BUS1_INTPRIO {
            display       "Interrupt priority of the SPI bus 1 ISR"
            flavor        data
            legal_values  0 to 15
            default_value 13
            description "
                This option specifies the interrupt priority of the ISR of
                the SPI bus 1 interrupt in the VIC. Slot 0 has the highest
                priority and slot 15 the lowest."
        }
    }

    cdl_component CYGPKG_DEVS_SPI_MICROBLAZE_OPTIONS {
        display "SPI build options"
        flavor  none
        no_define
    }

    cdl_option CYGPKG_DEVS_SPI_MICROBLAZE_TESTS {
        display         "SPI tests"
        flavor          data
        no_define
        calculated      { "tests/m25p05" }
        #tests/eth_test tests/spi 
#        default value {"tests/spi"}
    } 
}

# EOF spi_microblaze.cdl
