# ====================================================================
#
#      hal_microblaze_generic.cdl
#
#      Generic HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Michal Pfeifer
# Original data:  PowerPC
# Contributors:   gthomas
# Date:           1999-11-02
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_MICROBLAZE_GENERIC {
    display       "Platform generic support"
    include_dir   cyg/hal
    parent        CYGPKG_HAL_MICROBLAZE
    description   "
        Generic support."

    compile       plf_io.c hal_diag.c hal_aux.c platform.S \
                  src/xbasic_types.c src/xil_assert.c src/xil_io.c \
                  src/xintc.c src/xintc_g.c src/xintc_intr.c src/xintc_l.c src/xintc_options.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
# For now, until RedBoot is working
#    implements    CYGINT_HAL_USE_ROM_MONITOR_UNSUPPORTED


    cdl_option CYGNUM_HAL_UARTLITE {
        display       "Serial port of UART Lite"
        default_value 1
        active_if     { MON_UARTLITE_0 == 1 }
        compile       src/xuartlite_g.c src/xuartlite_intr.c \
            src/xuartlite_stats.c src/xuartlite.c src/xuartlite_l.c \
            src/xuartlite_selftest.c src/xuartlite_sinit.c
    }

    cdl_option CYGNUM_HAL_UART16550 {
        display       "Serial port of UART 16550"
        active_if     { MON_UART16550_0 == 1 }
        default_value 1
        compile       src/xuartns550_g.c src/xuartns550_intr.c \
            src/xuartns550_options.c  src/xuartns550_stats.c src/xuartns550.c src/xuartns550_l.c \
            src/xuartns550_selftest.c src/xuartns550_format.c src/xuartns550_sinit.c
    }

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_microblaze_platform.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLF_IO_H   <cyg/hal/plf_io.h>"
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM" "ROM" "ROMRAM"}
        default_value {"RAM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
           This option is used to control where the application program will
           run, either from RAM or ROM (flash) memory.  ROM based applications
           must be self contained, while RAM applications will typically assume
           the existence of a debug environment, such as GDB stubs."
    }

   cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
       display      "Number of communication channels on the board"
       flavor       data
       calculated   1
   }

   cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
       display          "Debug serial port"
       active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
       flavor data
       legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
       default_value    0
       description      "
           The board has only one serial port. This option
           chooses which port will be used to connect to a host
           running GDB."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
        display          "Diagnostic serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           The board has only one serial port.  This option
           chooses which port will be used for diagnostic output."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Baud rate for the HAL diagnostic port"
        flavor        data
        legal_values  { 50 75 110 "134_5" 150 200 300 600 1200 1800 2400 3600
                      4800 7200 9600 14400 19200 38400 57600 115200 230400
        }
        default_value 115200
        description   "
            This option specifies the default baud rate (speed) for the 
            HAL diagnostic port."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        description   "
            Period is busclock/100."
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            default_value 1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            default_value    { (MON_SYSTEM_CLK / 100) }
        }
        cdl_option CYGHWR_HAL_RTC_USE_AUTO_RESET {
            display       "Real-time clock timer use autoreset"
            flavor        bool
            default_value 1
            description   "
                This is best for precise time counting. If is autoreset true
                hal_clock_reset function do nothing if timer is running."
        }
    }
    
    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "microblazeel-unknown-linux-gnu" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
# -fvtable-gc -Woverloaded-virtual -Wstrict-prototypes    not supported in gcc
            default_value { CYGBLD_GLOBAL_WARNFLAGS . "-D__LITTLE_ENDIAN__ -fmessage-length=0 -mlittle-endian -mxl-barrel-shift -mno-xl-soft-mul \
				-g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -I. -I$(PREFIX)/include/cyg/hal/ " }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-fmessage-length=0 -mlittle-endian -mxl-barrel-shift -mno-xl-soft-mul -g -nostdlib -Wl,--gc-sections -Wl,-static" }
#            default_value { "-msoft-float -g -nostdlib" }
#            default_value { "-mcpu=v8.10.a -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the platform CDL takes care of creating
                an S-Record data file suitable for programming using
                the board's EPPC-Bug firmware monitor."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O srec --change-address=0x02000000 $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

#    cdl_component CYGPKG_HAL_MICROBLAZE_SPARTAN3ESK_OPTIONS {
#        display "SPARTAN3ESK build options"
#        flavor  none
#        description   "
#            Package specific build options including control over
#            compiler flags used only in building this package,
#            and details of which tests are built."
#    
#    
#        cdl_option CYGPKG_HAL_MICROBLAZE_SPARTAN3ESK_CFLAGS_ADD {
#            display "Additional compiler flags"
#            flavor  data
#            no_define
#            default_value { "" }
#            description   "
#                This option modifies the set of compiler flags for
#                building HAL. These flags are used in addition
#                to the set of global flags."
#        }
#    
#        cdl_option CYGPKG_HAL_MICROBLAZE_SPARTAN3ESK_CFLAGS_REMOVE {
#            display "Suppressed compiler flags"
#            flavor  data
#            no_define
#            default_value { "" }
#            description   "
#                This option modifies the set of compiler flags for
#                building HAL. These flags are removed from
#                the set of global flags if present."
#        }
#    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "microblaze_generic_ram" :
                                                "microblaze_generic_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_microblaze_generic_ram.ldi>" :
                                                    "<pkgconf/mlt_microblaze_generic_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_microblaze_generic_ram.h>" :
                                                    "<pkgconf/mlt_microblaze_generic_rom.h>" }
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" || CYG_HAL_STARTUP == "ROMRAM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

#        cdl_option CYGSEM_REDBOOT_PLF_LINUX_BOOT {
#            active_if      CYGBLD_BUILD_REDBOOT_WITH_EXEC
#            display        "Support booting Linux via RedBoot"
#            flavor         bool
#            default_value  1
#            description    "
#               This option enables RedBoot to support booting of a Linux kernel."
#
#            compile plf_redboot_linux_exec.c
#        }

        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 0
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to a binary image suitable for ROM programming."

#            compile -library=libextras.a redboot_cmds.c
 
            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img) 
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }
    }
}
