# ====================================================================
#
#      flash_at91eefc.cdl
#
#      FLASH programming for the Enhanced Embedded Flash Controller
#
# ====================================================================
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):
# Original data:
# Contributors:
# Date:
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_AT91EEFC {
    display      "AT91 EEFC FLASH memory support"

    parent       CYGPKG_IO_FLASH
    active_if    CYGPKG_IO_FLASH

    implements   CYGHWR_IO_FLASH_DEVICE

    include_dir  cyg/io

    description   "FLASH memory device support for AT91 EEFC"
    compile       at91eefc_flash.c
}
