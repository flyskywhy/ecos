# ====================================================================
#
#      devs_flash_at91sam9x25ek.cdl
#
#      FLASH memory - Hardware support NAND
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Denis Mikhayevich <denis.mikhayevich@axonim.by>
# Contributors:   
# Date:           2011-08-30
# Description:    FLASH drivers for NAND devices.
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_AT91SAN9X25EK { 
    display       "AT91SAN9X25EK NAND FLASH memory support" 
    description   "NAND FLASH memory device support for AT91SAN9X25EK" 
 
    include_dir   cyg/io 
 
    parent        CYGPKG_IO_FLASH 
    active_if     CYGPKG_IO_FLASH 
 
	define_proc { 
        puts $::cdl_system_header "#define CYGDAT_DEVS_FLASH_NAND_PLF_INL <cyg/io/devs_flash_at91sam9x25ek.inl>" 
    } 
 
   cdl_interface CYGINT_DEVS_FLASH_NAND_REQUIRED { 
       display   "NAND FLASH driver required" 
   } 
 
   implements    CYGINT_DEVS_FLASH_NAND_REQUIRED 
   implements    CYGHWR_IO_FLASH_DEVICE 
   implements	 CYGHWR_IO_FLASH_DEVICE_LEGACY
   implements    CYGHWR_IO_FLASH_INDIRECT_READS
} 

# EOF devs_flash_at91sam9x25ek.cdl